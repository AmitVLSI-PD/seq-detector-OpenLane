VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO seq_detector_mealy
  CLASS BLOCK ;
  FOREIGN seq_detector_mealy ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 19.115 10.640 20.715 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.310 10.640 42.910 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.505 10.640 65.105 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.700 10.640 87.300 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 22.900 94.540 24.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.940 94.540 43.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 60.980 94.540 62.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.020 94.540 81.620 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.600 94.540 21.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.640 94.540 40.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 57.680 94.540 59.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.720 94.540 78.320 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END clk
  PIN din
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END din
  PIN dout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.040 100.000 51.640 ;
    END
  END dout
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END reset
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 94.300 87.280 ;
      LAYER met2 ;
        RECT 15.845 4.280 92.830 87.225 ;
        RECT 15.845 4.000 48.110 4.280 ;
        RECT 48.950 4.000 92.830 4.280 ;
      LAYER met3 ;
        RECT 4.000 52.040 96.000 87.205 ;
        RECT 4.000 50.640 95.600 52.040 ;
        RECT 4.000 48.640 96.000 50.640 ;
        RECT 4.400 47.240 95.600 48.640 ;
        RECT 4.000 10.715 96.000 47.240 ;
  END
END seq_detector_mealy
END LIBRARY

