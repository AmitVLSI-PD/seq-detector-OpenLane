magic
tech sky130A
magscale 1 2
timestamp 1746547908
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 1104 2128 18860 17456
<< metal2 >>
rect 9678 0 9734 800
<< obsm2 >>
rect 3169 856 18566 17445
rect 3169 800 9622 856
rect 9790 800 18566 856
<< metal3 >>
rect 19200 10208 20000 10328
rect 0 9528 800 9648
rect 19200 9528 20000 9648
<< obsm3 >>
rect 800 10408 19200 17441
rect 800 10128 19120 10408
rect 800 9728 19200 10128
rect 880 9448 19120 9728
rect 800 2143 19200 9448
<< metal4 >>
rect 3163 2128 3483 17456
rect 3823 2128 4143 17456
rect 7602 2128 7922 17456
rect 8262 2128 8582 17456
rect 12041 2128 12361 17456
rect 12701 2128 13021 17456
rect 16480 2128 16800 17456
rect 17140 2128 17460 17456
<< metal5 >>
rect 1056 16004 18908 16324
rect 1056 15344 18908 15664
rect 1056 12196 18908 12516
rect 1056 11536 18908 11856
rect 1056 8388 18908 8708
rect 1056 7728 18908 8048
rect 1056 4580 18908 4900
rect 1056 3920 18908 4240
<< labels >>
rlabel metal4 s 3823 2128 4143 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8262 2128 8582 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12701 2128 13021 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17140 2128 17460 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4580 18908 4900 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8388 18908 8708 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12196 18908 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16004 18908 16324 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3163 2128 3483 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3920 18908 4240 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7728 18908 8048 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11536 18908 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15344 18908 15664 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 9528 800 9648 6 clk
port 3 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 din
port 4 nsew signal input
rlabel metal3 s 19200 10208 20000 10328 6 dout
port 5 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 reset
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 291936
string GDS_FILE /openlane/designs/seq_detector/runs/RUN_2025.05.06_16.09.42/results/signoff/seq_detector_mealy.magic.gds
string GDS_START 87230
<< end >>

